library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.IDecode_const.all;

package rom is

constant ROM_SIZE : integer := 22;
TYPE ROM is array(0 to ROM_SIZE - 1) of std_logic_vector(31 downto 0);

constant boot_rom : ROM := (
X"00000000",
F_LUI  &"00000"&"11111"&X"0000",
F_ADDIU&"11111"&"00000"&X"0007",
F_ADDIU&"11111"&"00001"&X"0000",
F_MFC0 &"00100"&"00000"&"00001"&"00000"&"000000",
F_LUI  &"00000"&"00000"&X"a000",
F_ADDIU&"11111"&"00001"&X"000a",
F_MFC0 &"00100"&"00000"&"00001"&"00000"&"000000",
F_ADDIU&"11111"&"00000"&X"0002",
F_ADDIU&"11111"&"00001"&X"0003",
F_MFC0 &"00100"&"00000"&"00001"&"00000"&"000000",
F_ADDIU&"11111"&"00000"&X"0002",
F_ADDIU&"11111"&"00001"&X"0002",
F_MFC0 &"00100"&"00000"&"00001"&"00000"&"000000",
F_TLBWI&"10000"&"00000"&"00000"&"00000"&"000010",
F_ADDIU&"11111"&"00000"&X"F0F0",
F_LUI  &"00000"&"00001"&X"a000",--92
F_SW   &"00001"&"00000"&X"0000",--93
F_LW   &"00001"&"00010"&X"0000",--94
F_MFC0 &"00000"&"00000"&"00001"&"00000"&"000000",--95
F_BNE  &"00000"&"00001"&X"ffec",
X"00000000"
    );

end rom;


